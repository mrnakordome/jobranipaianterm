library verilog;
use verilog.vl_types.all;
entity TBQ7 is
end TBQ7;
